library IEEE;
use IEEE.STD_LOGIC_1164.ALL;


entity XNOR_GATE is 
port
(

INPUT_A ,INPUT_B : IN STD_LOGIC;
OUTPUT : OUT STD_LOGIC

);

end XNOR_GATE;

Architecture behavioral of XNOR_GATE is begin

OUTPUT<= INPUT_A XNOR INPUT_B;

end behavioral;

